/*
 * gemm_layer design including complex dsp definition
*/

`define complex_dsp

`include "./generic_circuits/gemm_layer.v"
