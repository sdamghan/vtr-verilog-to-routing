/*
 * eltwise_layer design including complex dsp definition
*/

`define complex_dsp

`include "./generic_circuits/eltwise_layer.v"
