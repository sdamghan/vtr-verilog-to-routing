module logical_left_shift_const (
				input   [71:0]	   unsigned_a,
                                output [63:0] unsigned_left_shift
                           );

    assign    unsigned_left_shift  =   unsigned_a << 65;

endmodule
