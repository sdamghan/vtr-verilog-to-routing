module signed_arithmetic_left_shift_variable (
				input [15:0]	shift,
				input  signed  [71:0]	   signed_a,
                                output signed [63:0] signed_left_shift
                           );

    assign    signed_left_shift  =   signed_a <<< shift[8:0];

endmodule
