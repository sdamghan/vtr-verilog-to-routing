/*
 * attention_layer design including complex dsp definition
*/

`define complex_dsp

`include "./generic_circuits/attention_layer.v"
