/*
 * robot_rl design including complex dsp definition
*/

`define complex_dsp

`include "./generic_circuits/robot_rl.v"
