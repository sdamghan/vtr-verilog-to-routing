/*
 * softmax design including complex dsp definition
*/

`define complex_dsp

`include "./generic_circuits/softmax.v"
